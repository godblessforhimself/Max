library verilog;
use verilog.vl_types.all;
entity vga640480_vlg_vec_tst is
end vga640480_vlg_vec_tst;
